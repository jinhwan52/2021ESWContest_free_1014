// nios2.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module nios2 (
		output wire        adc_ltc2308_0_conduit_end_CONVST,             //             adc_ltc2308_0_conduit_end.CONVST
		output wire        adc_ltc2308_0_conduit_end_SCK,                //                                      .SCK
		output wire        adc_ltc2308_0_conduit_end_SDI,                //                                      .SDI
		input  wire        adc_ltc2308_0_conduit_end_SDO,                //                                      .SDO
		input  wire [4:0]  bridge_0_external_interface_address,          //           bridge_0_external_interface.address
		input  wire [1:0]  bridge_0_external_interface_byte_enable,      //                                      .byte_enable
		input  wire        bridge_0_external_interface_read,             //                                      .read
		input  wire        bridge_0_external_interface_write,            //                                      .write
		input  wire [15:0] bridge_0_external_interface_write_data,       //                                      .write_data
		output wire        bridge_0_external_interface_acknowledge,      //                                      .acknowledge
		output wire [15:0] bridge_0_external_interface_read_data,        //                                      .read_data
		input  wire        clk_clk,                                      //                                   clk.clk
		input  wire        clock_bridge_0_in_clk_clk,                    //                 clock_bridge_0_in_clk.clk
		output wire        clock_bridge_100_out_clk_clk,                 //              clock_bridge_100_out_clk.clk
		output wire        clock_bridge_65_out_clk_clk,                  //               clock_bridge_65_out_clk.clk
		output wire [31:0] command_from_hps_external_connection_export,  //  command_from_hps_external_connection.export
		output wire [31:0] electrode_voltage_external_connection_export, // electrode_voltage_external_connection.export
		input  wire        fifo_fpga_to_hps_clk_in_clk,                  //               fifo_fpga_to_hps_clk_in.clk
		input  wire [31:0] fifo_fpga_to_hps_in_writedata,                //                   fifo_fpga_to_hps_in.writedata
		input  wire        fifo_fpga_to_hps_in_write,                    //                                      .write
		input  wire [2:0]  fifo_fpga_to_hps_in_csr_address,              //               fifo_fpga_to_hps_in_csr.address
		input  wire        fifo_fpga_to_hps_in_csr_read,                 //                                      .read
		input  wire [31:0] fifo_fpga_to_hps_in_csr_writedata,            //                                      .writedata
		input  wire        fifo_fpga_to_hps_in_csr_write,                //                                      .write
		output wire [31:0] fifo_fpga_to_hps_in_csr_readdata,             //                                      .readdata
		input  wire        fifo_fpga_to_hps_reset_in_reset_n,            //             fifo_fpga_to_hps_reset_in.reset_n
		input  wire        fifo_hps_to_fpga_clk_out_clk,                 //              fifo_hps_to_fpga_clk_out.clk
		output wire [31:0] fifo_hps_to_fpga_out_readdata,                //                  fifo_hps_to_fpga_out.readdata
		input  wire        fifo_hps_to_fpga_out_read,                    //                                      .read
		input  wire [2:0]  fifo_hps_to_fpga_out_csr_address,             //              fifo_hps_to_fpga_out_csr.address
		input  wire        fifo_hps_to_fpga_out_csr_read,                //                                      .read
		input  wire [31:0] fifo_hps_to_fpga_out_csr_writedata,           //                                      .writedata
		input  wire        fifo_hps_to_fpga_out_csr_write,               //                                      .write
		output wire [31:0] fifo_hps_to_fpga_out_csr_readdata,            //                                      .readdata
		input  wire        fifo_hps_to_fpga_reset_out_reset_n,           //            fifo_hps_to_fpga_reset_out.reset_n
		input  wire [7:0]  finish_fdtd_external_connection_export,       //       finish_fdtd_external_connection.export
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,              //                                hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,                //                                      .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,                //                                      .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,                //                                      .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,                //                                      .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,                //                                      .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,                //                                      .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,                 //                                      .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,              //                                      .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,              //                                      .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,              //                                      .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,                //                                      .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,                //                                      .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,                //                                      .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,                  //                                      .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,                  //                                      .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,                  //                                      .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,                  //                                      .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,                  //                                      .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,                  //                                      .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,                  //                                      .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,                   //                                      .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,                   //                                      .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,                  //                                      .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,                   //                                      .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,                   //                                      .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,                   //                                      .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,                   //                                      .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,                   //                                      .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,                   //                                      .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,                   //                                      .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,                   //                                      .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,                   //                                      .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,                   //                                      .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,                  //                                      .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,                  //                                      .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,                  //                                      .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,                  //                                      .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,                 //                                      .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,                //                                      .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,                //                                      .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,                 //                                      .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,                  //                                      .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,                  //                                      .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,                  //                                      .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,                  //                                      .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,                  //                                      .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,                  //                                      .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,               //                                      .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,               //                                      .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,               //                                      .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,               //                                      .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,               //                                      .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,               //                                      .hps_io_gpio_inst_GPIO61
		output wire [7:0]  hw_reset_external_connection_export,          //          hw_reset_external_connection.export
		output wire [15:0] iteration_number_external_connection_export,  //  iteration_number_external_connection.export
		output wire [14:0] memory_mem_a,                                 //                                memory.mem_a
		output wire [2:0]  memory_mem_ba,                                //                                      .mem_ba
		output wire        memory_mem_ck,                                //                                      .mem_ck
		output wire        memory_mem_ck_n,                              //                                      .mem_ck_n
		output wire        memory_mem_cke,                               //                                      .mem_cke
		output wire        memory_mem_cs_n,                              //                                      .mem_cs_n
		output wire        memory_mem_ras_n,                             //                                      .mem_ras_n
		output wire        memory_mem_cas_n,                             //                                      .mem_cas_n
		output wire        memory_mem_we_n,                              //                                      .mem_we_n
		output wire        memory_mem_reset_n,                           //                                      .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                                //                                      .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                               //                                      .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                             //                                      .mem_dqs_n
		output wire        memory_mem_odt,                               //                                      .mem_odt
		output wire [3:0]  memory_mem_dm,                                //                                      .mem_dm
		input  wire        memory_oct_rzqin,                             //                                      .oct_rzqin
		input  wire [15:0] module_csr_external_connection_export,        //        module_csr_external_connection.export
		input  wire [31:0] number32_export,                              //                              number32.export
		input  wire [15:0] o_pw_forward_external_connection_export,      //      o_pw_forward_external_connection.export
		input  wire [15:0] o_pw_reversed_external_connection_export,     //     o_pw_reversed_external_connection.export
		input  wire [15:0] o_temperature2_external_connection_export,    //    o_temperature2_external_connection.export
		input  wire [15:0] o_temperature_external_connection_export,     //     o_temperature_external_connection.export
		input  wire        onchip_ram1_reset1_reset,                     //                    onchip_ram1_reset1.reset
		input  wire        onchip_ram1_reset1_reset_req,                 //                                      .reset_req
		input  wire [6:0]  onchip_ram1_s1_address,                       //                        onchip_ram1_s1.address
		input  wire        onchip_ram1_s1_clken,                         //                                      .clken
		input  wire        onchip_ram1_s1_chipselect,                    //                                      .chipselect
		input  wire        onchip_ram1_s1_write,                         //                                      .write
		output wire [15:0] onchip_ram1_s1_readdata,                      //                                      .readdata
		input  wire [15:0] onchip_ram1_s1_writedata,                     //                                      .writedata
		input  wire [1:0]  onchip_ram1_s1_byteenable,                    //                                      .byteenable
		input  wire        onchip_ram2_reset1_reset,                     //                    onchip_ram2_reset1.reset
		input  wire        onchip_ram2_reset1_reset_req,                 //                                      .reset_req
		input  wire [6:0]  onchip_ram2_s1_address,                       //                        onchip_ram2_s1.address
		input  wire        onchip_ram2_s1_clken,                         //                                      .clken
		input  wire        onchip_ram2_s1_chipselect,                    //                                      .chipselect
		input  wire        onchip_ram2_s1_write,                         //                                      .write
		output wire [15:0] onchip_ram2_s1_readdata,                      //                                      .readdata
		input  wire [15:0] onchip_ram2_s1_writedata,                     //                                      .writedata
		input  wire [1:0]  onchip_ram2_s1_byteenable,                    //                                      .byteenable
		output wire        pll_adc_locked_export,                        //                        pll_adc_locked.export
		output wire [7:0]  power_unlock_external_connection_export,      //      power_unlock_external_connection.export
		input  wire        reset_reset,                                  //                                 reset.reset
		output wire        rf_on_off_external_connection_export,         //         rf_on_off_external_connection.export
		output wire        sdram_clk_clk,                                //                             sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                              //                            sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                //                                      .ba
		output wire        sdram_wire_cas_n,                             //                                      .cas_n
		output wire        sdram_wire_cke,                               //                                      .cke
		output wire        sdram_wire_cs_n,                              //                                      .cs_n
		inout  wire [15:0] sdram_wire_dq,                                //                                      .dq
		output wire [1:0]  sdram_wire_dqm,                               //                                      .dqm
		output wire        sdram_wire_ras_n,                             //                                      .ras_n
		output wire        sdram_wire_we_n,                              //                                      .we_n
		output wire [19:0] sp_external_connection_export,                //                sp_external_connection.export
		input  wire [9:0]  sw_external_connection_export,                //                sw_external_connection.export
		output wire        thermocouples_sel_external_connection_export, // thermocouples_sel_external_connection.export
		output wire        vga_out_CLK,                                  //                               vga_out.CLK
		output wire        vga_out_HS,                                   //                                      .HS
		output wire        vga_out_VS,                                   //                                      .VS
		output wire        vga_out_BLANK,                                //                                      .BLANK
		output wire        vga_out_SYNC,                                 //                                      .SYNC
		output wire [7:0]  vga_out_R,                                    //                                      .R
		output wire [7:0]  vga_out_G,                                    //                                      .G
		output wire [7:0]  vga_out_B,                                    //                                      .B
		input  wire        vga_ref_reset_reset,                          //                         vga_ref_reset.reset
		input  wire        video_ref_clk_clk                             //                         video_ref_clk.clk
	);

	wire          pll_adc_outclk0_clk;                                            // pll_adc:outclk_0 -> temperature_adc:adc_clk
	wire   [15:0] bridge_fpga_tempadc_avalon_master_readdata;                     // mm_interconnect_0:bridge_FPGA_tempADC_avalon_master_readdata -> bridge_FPGA_tempADC:avalon_readdata
	wire          bridge_fpga_tempadc_avalon_master_waitrequest;                  // mm_interconnect_0:bridge_FPGA_tempADC_avalon_master_waitrequest -> bridge_FPGA_tempADC:avalon_waitrequest
	wire    [1:0] bridge_fpga_tempadc_avalon_master_byteenable;                   // bridge_FPGA_tempADC:avalon_byteenable -> mm_interconnect_0:bridge_FPGA_tempADC_avalon_master_byteenable
	wire          bridge_fpga_tempadc_avalon_master_read;                         // bridge_FPGA_tempADC:avalon_read -> mm_interconnect_0:bridge_FPGA_tempADC_avalon_master_read
	wire    [4:0] bridge_fpga_tempadc_avalon_master_address;                      // bridge_FPGA_tempADC:avalon_address -> mm_interconnect_0:bridge_FPGA_tempADC_avalon_master_address
	wire          bridge_fpga_tempadc_avalon_master_write;                        // bridge_FPGA_tempADC:avalon_write -> mm_interconnect_0:bridge_FPGA_tempADC_avalon_master_write
	wire   [15:0] bridge_fpga_tempadc_avalon_master_writedata;                    // bridge_FPGA_tempADC:avalon_writedata -> mm_interconnect_0:bridge_FPGA_tempADC_avalon_master_writedata
	wire          mm_interconnect_0_temperature_adc_slave_chipselect;             // mm_interconnect_0:temperature_adc_slave_chipselect -> temperature_adc:slave_chipselect_n
	wire   [15:0] mm_interconnect_0_temperature_adc_slave_readdata;               // temperature_adc:slave_readdata -> mm_interconnect_0:temperature_adc_slave_readdata
	wire    [0:0] mm_interconnect_0_temperature_adc_slave_address;                // mm_interconnect_0:temperature_adc_slave_address -> temperature_adc:slave_addr
	wire          mm_interconnect_0_temperature_adc_slave_read;                   // mm_interconnect_0:temperature_adc_slave_read -> temperature_adc:slave_read_n
	wire          mm_interconnect_0_temperature_adc_slave_write;                  // mm_interconnect_0:temperature_adc_slave_write -> temperature_adc:slave_wrtie_n
	wire   [15:0] mm_interconnect_0_temperature_adc_slave_writedata;              // mm_interconnect_0:temperature_adc_slave_writedata -> temperature_adc:slave_wriredata
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                   // hps_0:h2f_AWBURST -> mm_interconnect_1:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                     // hps_0:h2f_ARLEN -> mm_interconnect_1:hps_0_h2f_axi_master_arlen
	wire   [15:0] hps_0_h2f_axi_master_wstrb;                                     // hps_0:h2f_WSTRB -> mm_interconnect_1:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                                    // mm_interconnect_1:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                       // mm_interconnect_1:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                                    // hps_0:h2f_RREADY -> mm_interconnect_1:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                     // hps_0:h2f_AWLEN -> mm_interconnect_1:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                       // hps_0:h2f_WID -> mm_interconnect_1:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                   // hps_0:h2f_ARCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                                    // hps_0:h2f_WVALID -> mm_interconnect_1:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                    // hps_0:h2f_ARADDR -> mm_interconnect_1:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                    // hps_0:h2f_ARPROT -> mm_interconnect_1:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                    // hps_0:h2f_AWPROT -> mm_interconnect_1:hps_0_h2f_axi_master_awprot
	wire  [127:0] hps_0_h2f_axi_master_wdata;                                     // hps_0:h2f_WDATA -> mm_interconnect_1:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                                   // hps_0:h2f_ARVALID -> mm_interconnect_1:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                   // hps_0:h2f_AWCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                                      // hps_0:h2f_ARID -> mm_interconnect_1:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                    // hps_0:h2f_ARLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                    // hps_0:h2f_AWLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                    // hps_0:h2f_AWADDR -> mm_interconnect_1:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                     // mm_interconnect_1:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                                   // mm_interconnect_1:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [127:0] hps_0_h2f_axi_master_rdata;                                     // mm_interconnect_1:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                                   // mm_interconnect_1:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                   // hps_0:h2f_ARBURST -> mm_interconnect_1:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                    // hps_0:h2f_ARSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                                    // hps_0:h2f_BREADY -> mm_interconnect_1:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                                     // mm_interconnect_1:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                                     // hps_0:h2f_WLAST -> mm_interconnect_1:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                     // mm_interconnect_1:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                                      // hps_0:h2f_AWID -> mm_interconnect_1:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                       // mm_interconnect_1:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                                    // mm_interconnect_1:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                    // hps_0:h2f_AWSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                                   // hps_0:h2f_AWVALID -> mm_interconnect_1:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                                    // mm_interconnect_1:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire          vga_subsystem_pixel_dma_master_waitrequest;                     // mm_interconnect_1:VGA_subsystem_pixel_dma_master_waitrequest -> VGA_subsystem:pixel_dma_master_waitrequest
	wire   [15:0] vga_subsystem_pixel_dma_master_readdata;                        // mm_interconnect_1:VGA_subsystem_pixel_dma_master_readdata -> VGA_subsystem:pixel_dma_master_readdata
	wire   [31:0] vga_subsystem_pixel_dma_master_address;                         // VGA_subsystem:pixel_dma_master_address -> mm_interconnect_1:VGA_subsystem_pixel_dma_master_address
	wire          vga_subsystem_pixel_dma_master_read;                            // VGA_subsystem:pixel_dma_master_read -> mm_interconnect_1:VGA_subsystem_pixel_dma_master_read
	wire          vga_subsystem_pixel_dma_master_readdatavalid;                   // mm_interconnect_1:VGA_subsystem_pixel_dma_master_readdatavalid -> VGA_subsystem:pixel_dma_master_readdatavalid
	wire          vga_subsystem_pixel_dma_master_lock;                            // VGA_subsystem:pixel_dma_master_lock -> mm_interconnect_1:VGA_subsystem_pixel_dma_master_lock
	wire          mm_interconnect_1_vga_subsystem_char_buffer_slave_chipselect;   // mm_interconnect_1:VGA_subsystem_char_buffer_slave_chipselect -> VGA_subsystem:char_buffer_slave_chipselect
	wire    [7:0] mm_interconnect_1_vga_subsystem_char_buffer_slave_readdata;     // VGA_subsystem:char_buffer_slave_readdata -> mm_interconnect_1:VGA_subsystem_char_buffer_slave_readdata
	wire          mm_interconnect_1_vga_subsystem_char_buffer_slave_waitrequest;  // VGA_subsystem:char_buffer_slave_waitrequest -> mm_interconnect_1:VGA_subsystem_char_buffer_slave_waitrequest
	wire   [12:0] mm_interconnect_1_vga_subsystem_char_buffer_slave_address;      // mm_interconnect_1:VGA_subsystem_char_buffer_slave_address -> VGA_subsystem:char_buffer_slave_address
	wire          mm_interconnect_1_vga_subsystem_char_buffer_slave_read;         // mm_interconnect_1:VGA_subsystem_char_buffer_slave_read -> VGA_subsystem:char_buffer_slave_read
	wire    [0:0] mm_interconnect_1_vga_subsystem_char_buffer_slave_byteenable;   // mm_interconnect_1:VGA_subsystem_char_buffer_slave_byteenable -> VGA_subsystem:char_buffer_slave_byteenable
	wire          mm_interconnect_1_vga_subsystem_char_buffer_slave_write;        // mm_interconnect_1:VGA_subsystem_char_buffer_slave_write -> VGA_subsystem:char_buffer_slave_write
	wire    [7:0] mm_interconnect_1_vga_subsystem_char_buffer_slave_writedata;    // mm_interconnect_1:VGA_subsystem_char_buffer_slave_writedata -> VGA_subsystem:char_buffer_slave_writedata
	wire          mm_interconnect_1_fifo_hps_to_fpga_in_write;                    // mm_interconnect_1:fifo_HPS_to_FPGA_in_write -> fifo_HPS_to_FPGA:avalonmm_write_slave_write
	wire   [31:0] mm_interconnect_1_fifo_hps_to_fpga_in_writedata;                // mm_interconnect_1:fifo_HPS_to_FPGA_in_writedata -> fifo_HPS_to_FPGA:avalonmm_write_slave_writedata
	wire   [31:0] mm_interconnect_1_fifo_fpga_to_hps_out_readdata;                // fifo_FPGA_to_HPS:avalonmm_read_slave_readdata -> mm_interconnect_1:fifo_FPGA_to_HPS_out_readdata
	wire          mm_interconnect_1_fifo_fpga_to_hps_out_read;                    // mm_interconnect_1:fifo_FPGA_to_HPS_out_read -> fifo_FPGA_to_HPS:avalonmm_read_slave_read
	wire          mm_interconnect_1_sdram_s1_chipselect;                          // mm_interconnect_1:sdram_s1_chipselect -> sdram:az_cs
	wire   [15:0] mm_interconnect_1_sdram_s1_readdata;                            // sdram:za_data -> mm_interconnect_1:sdram_s1_readdata
	wire          mm_interconnect_1_sdram_s1_waitrequest;                         // sdram:za_waitrequest -> mm_interconnect_1:sdram_s1_waitrequest
	wire   [24:0] mm_interconnect_1_sdram_s1_address;                             // mm_interconnect_1:sdram_s1_address -> sdram:az_addr
	wire          mm_interconnect_1_sdram_s1_read;                                // mm_interconnect_1:sdram_s1_read -> sdram:az_rd_n
	wire    [1:0] mm_interconnect_1_sdram_s1_byteenable;                          // mm_interconnect_1:sdram_s1_byteenable -> sdram:az_be_n
	wire          mm_interconnect_1_sdram_s1_readdatavalid;                       // sdram:za_valid -> mm_interconnect_1:sdram_s1_readdatavalid
	wire          mm_interconnect_1_sdram_s1_write;                               // mm_interconnect_1:sdram_s1_write -> sdram:az_wr_n
	wire   [15:0] mm_interconnect_1_sdram_s1_writedata;                           // mm_interconnect_1:sdram_s1_writedata -> sdram:az_data
	wire          mm_interconnect_1_onchip_ram1_s2_chipselect;                    // mm_interconnect_1:onchip_ram1_s2_chipselect -> onchip_ram1:chipselect2
	wire   [15:0] mm_interconnect_1_onchip_ram1_s2_readdata;                      // onchip_ram1:readdata2 -> mm_interconnect_1:onchip_ram1_s2_readdata
	wire    [6:0] mm_interconnect_1_onchip_ram1_s2_address;                       // mm_interconnect_1:onchip_ram1_s2_address -> onchip_ram1:address2
	wire    [1:0] mm_interconnect_1_onchip_ram1_s2_byteenable;                    // mm_interconnect_1:onchip_ram1_s2_byteenable -> onchip_ram1:byteenable2
	wire          mm_interconnect_1_onchip_ram1_s2_write;                         // mm_interconnect_1:onchip_ram1_s2_write -> onchip_ram1:write2
	wire   [15:0] mm_interconnect_1_onchip_ram1_s2_writedata;                     // mm_interconnect_1:onchip_ram1_s2_writedata -> onchip_ram1:writedata2
	wire          mm_interconnect_1_onchip_ram1_s2_clken;                         // mm_interconnect_1:onchip_ram1_s2_clken -> onchip_ram1:clken2
	wire          mm_interconnect_1_onchip_ram2_s2_chipselect;                    // mm_interconnect_1:onchip_ram2_s2_chipselect -> onchip_ram2:chipselect2
	wire   [15:0] mm_interconnect_1_onchip_ram2_s2_readdata;                      // onchip_ram2:readdata2 -> mm_interconnect_1:onchip_ram2_s2_readdata
	wire    [6:0] mm_interconnect_1_onchip_ram2_s2_address;                       // mm_interconnect_1:onchip_ram2_s2_address -> onchip_ram2:address2
	wire    [1:0] mm_interconnect_1_onchip_ram2_s2_byteenable;                    // mm_interconnect_1:onchip_ram2_s2_byteenable -> onchip_ram2:byteenable2
	wire          mm_interconnect_1_onchip_ram2_s2_write;                         // mm_interconnect_1:onchip_ram2_s2_write -> onchip_ram2:write2
	wire   [15:0] mm_interconnect_1_onchip_ram2_s2_writedata;                     // mm_interconnect_1:onchip_ram2_s2_writedata -> onchip_ram2:writedata2
	wire          mm_interconnect_1_onchip_ram2_s2_clken;                         // mm_interconnect_1:onchip_ram2_s2_clken -> onchip_ram2:clken2
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                                // hps_0:h2f_lw_AWBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                  // hps_0:h2f_lw_ARLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                  // hps_0:h2f_lw_WSTRB -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                                 // mm_interconnect_2:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                    // mm_interconnect_2:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                                 // hps_0:h2f_lw_RREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                  // hps_0:h2f_lw_AWLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                    // hps_0:h2f_lw_WID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                                // hps_0:h2f_lw_ARCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                                 // hps_0:h2f_lw_WVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                 // hps_0:h2f_lw_ARADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                 // hps_0:h2f_lw_ARPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                 // hps_0:h2f_lw_AWPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                  // hps_0:h2f_lw_WDATA -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                                // hps_0:h2f_lw_ARVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                                // hps_0:h2f_lw_AWCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                   // hps_0:h2f_lw_ARID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                 // hps_0:h2f_lw_ARLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                 // hps_0:h2f_lw_AWLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                 // hps_0:h2f_lw_AWADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                  // mm_interconnect_2:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                                // mm_interconnect_2:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                  // mm_interconnect_2:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                                // mm_interconnect_2:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                                // hps_0:h2f_lw_ARBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                 // hps_0:h2f_lw_ARSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                                 // hps_0:h2f_lw_BREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                                  // mm_interconnect_2:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                                  // hps_0:h2f_lw_WLAST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                  // mm_interconnect_2:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                   // hps_0:h2f_lw_AWID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                    // mm_interconnect_2:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                                 // mm_interconnect_2:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                 // hps_0:h2f_lw_AWSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                                // hps_0:h2f_lw_AWVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                                 // mm_interconnect_2:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire          mm_interconnect_2_vga_subsystem_char_control_slave_chipselect;  // mm_interconnect_2:VGA_subsystem_char_control_slave_chipselect -> VGA_subsystem:char_control_slave_chipselect
	wire   [31:0] mm_interconnect_2_vga_subsystem_char_control_slave_readdata;    // VGA_subsystem:char_control_slave_readdata -> mm_interconnect_2:VGA_subsystem_char_control_slave_readdata
	wire    [0:0] mm_interconnect_2_vga_subsystem_char_control_slave_address;     // mm_interconnect_2:VGA_subsystem_char_control_slave_address -> VGA_subsystem:char_control_slave_address
	wire          mm_interconnect_2_vga_subsystem_char_control_slave_read;        // mm_interconnect_2:VGA_subsystem_char_control_slave_read -> VGA_subsystem:char_control_slave_read
	wire    [3:0] mm_interconnect_2_vga_subsystem_char_control_slave_byteenable;  // mm_interconnect_2:VGA_subsystem_char_control_slave_byteenable -> VGA_subsystem:char_control_slave_byteenable
	wire          mm_interconnect_2_vga_subsystem_char_control_slave_write;       // mm_interconnect_2:VGA_subsystem_char_control_slave_write -> VGA_subsystem:char_control_slave_write
	wire   [31:0] mm_interconnect_2_vga_subsystem_char_control_slave_writedata;   // mm_interconnect_2:VGA_subsystem_char_control_slave_writedata -> VGA_subsystem:char_control_slave_writedata
	wire   [31:0] mm_interconnect_2_fifo_hps_to_fpga_in_csr_readdata;             // fifo_HPS_to_FPGA:wrclk_control_slave_readdata -> mm_interconnect_2:fifo_HPS_to_FPGA_in_csr_readdata
	wire    [2:0] mm_interconnect_2_fifo_hps_to_fpga_in_csr_address;              // mm_interconnect_2:fifo_HPS_to_FPGA_in_csr_address -> fifo_HPS_to_FPGA:wrclk_control_slave_address
	wire          mm_interconnect_2_fifo_hps_to_fpga_in_csr_read;                 // mm_interconnect_2:fifo_HPS_to_FPGA_in_csr_read -> fifo_HPS_to_FPGA:wrclk_control_slave_read
	wire          mm_interconnect_2_fifo_hps_to_fpga_in_csr_write;                // mm_interconnect_2:fifo_HPS_to_FPGA_in_csr_write -> fifo_HPS_to_FPGA:wrclk_control_slave_write
	wire   [31:0] mm_interconnect_2_fifo_hps_to_fpga_in_csr_writedata;            // mm_interconnect_2:fifo_HPS_to_FPGA_in_csr_writedata -> fifo_HPS_to_FPGA:wrclk_control_slave_writedata
	wire   [31:0] mm_interconnect_2_fifo_fpga_to_hps_out_csr_readdata;            // fifo_FPGA_to_HPS:rdclk_control_slave_readdata -> mm_interconnect_2:fifo_FPGA_to_HPS_out_csr_readdata
	wire    [2:0] mm_interconnect_2_fifo_fpga_to_hps_out_csr_address;             // mm_interconnect_2:fifo_FPGA_to_HPS_out_csr_address -> fifo_FPGA_to_HPS:rdclk_control_slave_address
	wire          mm_interconnect_2_fifo_fpga_to_hps_out_csr_read;                // mm_interconnect_2:fifo_FPGA_to_HPS_out_csr_read -> fifo_FPGA_to_HPS:rdclk_control_slave_read
	wire          mm_interconnect_2_fifo_fpga_to_hps_out_csr_write;               // mm_interconnect_2:fifo_FPGA_to_HPS_out_csr_write -> fifo_FPGA_to_HPS:rdclk_control_slave_write
	wire   [31:0] mm_interconnect_2_fifo_fpga_to_hps_out_csr_writedata;           // mm_interconnect_2:fifo_FPGA_to_HPS_out_csr_writedata -> fifo_FPGA_to_HPS:rdclk_control_slave_writedata
	wire   [31:0] mm_interconnect_2_sw_s1_readdata;                               // SW:readdata -> mm_interconnect_2:SW_s1_readdata
	wire    [1:0] mm_interconnect_2_sw_s1_address;                                // mm_interconnect_2:SW_s1_address -> SW:address
	wire   [31:0] mm_interconnect_2_number32_s1_readdata;                         // Number32:readdata -> mm_interconnect_2:Number32_s1_readdata
	wire    [1:0] mm_interconnect_2_number32_s1_address;                          // mm_interconnect_2:Number32_s1_address -> Number32:address
	wire   [31:0] mm_interconnect_2_o_temperature_s1_readdata;                    // O_temperature:readdata -> mm_interconnect_2:O_temperature_s1_readdata
	wire    [1:0] mm_interconnect_2_o_temperature_s1_address;                     // mm_interconnect_2:O_temperature_s1_address -> O_temperature:address
	wire   [31:0] mm_interconnect_2_o_pw_forward_s1_readdata;                     // O_pw_forward:readdata -> mm_interconnect_2:O_pw_forward_s1_readdata
	wire    [1:0] mm_interconnect_2_o_pw_forward_s1_address;                      // mm_interconnect_2:O_pw_forward_s1_address -> O_pw_forward:address
	wire   [31:0] mm_interconnect_2_o_pw_reversed_s1_readdata;                    // O_pw_reversed:readdata -> mm_interconnect_2:O_pw_reversed_s1_readdata
	wire    [1:0] mm_interconnect_2_o_pw_reversed_s1_address;                     // mm_interconnect_2:O_pw_reversed_s1_address -> O_pw_reversed:address
	wire   [31:0] mm_interconnect_2_o_temperature2_s1_readdata;                   // O_temperature2:readdata -> mm_interconnect_2:O_temperature2_s1_readdata
	wire    [1:0] mm_interconnect_2_o_temperature2_s1_address;                    // mm_interconnect_2:O_temperature2_s1_address -> O_temperature2:address
	wire          mm_interconnect_2_rf_on_off_s1_chipselect;                      // mm_interconnect_2:rf_on_off_s1_chipselect -> rf_on_off:chipselect
	wire   [31:0] mm_interconnect_2_rf_on_off_s1_readdata;                        // rf_on_off:readdata -> mm_interconnect_2:rf_on_off_s1_readdata
	wire    [1:0] mm_interconnect_2_rf_on_off_s1_address;                         // mm_interconnect_2:rf_on_off_s1_address -> rf_on_off:address
	wire          mm_interconnect_2_rf_on_off_s1_write;                           // mm_interconnect_2:rf_on_off_s1_write -> rf_on_off:write_n
	wire   [31:0] mm_interconnect_2_rf_on_off_s1_writedata;                       // mm_interconnect_2:rf_on_off_s1_writedata -> rf_on_off:writedata
	wire          mm_interconnect_2_command_from_hps_s1_chipselect;               // mm_interconnect_2:command_from_hps_s1_chipselect -> command_from_hps:chipselect
	wire   [31:0] mm_interconnect_2_command_from_hps_s1_readdata;                 // command_from_hps:readdata -> mm_interconnect_2:command_from_hps_s1_readdata
	wire    [1:0] mm_interconnect_2_command_from_hps_s1_address;                  // mm_interconnect_2:command_from_hps_s1_address -> command_from_hps:address
	wire          mm_interconnect_2_command_from_hps_s1_write;                    // mm_interconnect_2:command_from_hps_s1_write -> command_from_hps:write_n
	wire   [31:0] mm_interconnect_2_command_from_hps_s1_writedata;                // mm_interconnect_2:command_from_hps_s1_writedata -> command_from_hps:writedata
	wire          mm_interconnect_2_sp_s1_chipselect;                             // mm_interconnect_2:SP_s1_chipselect -> SP:chipselect
	wire   [31:0] mm_interconnect_2_sp_s1_readdata;                               // SP:readdata -> mm_interconnect_2:SP_s1_readdata
	wire    [1:0] mm_interconnect_2_sp_s1_address;                                // mm_interconnect_2:SP_s1_address -> SP:address
	wire          mm_interconnect_2_sp_s1_write;                                  // mm_interconnect_2:SP_s1_write -> SP:write_n
	wire   [31:0] mm_interconnect_2_sp_s1_writedata;                              // mm_interconnect_2:SP_s1_writedata -> SP:writedata
	wire          mm_interconnect_2_thermocouples_sel_s1_chipselect;              // mm_interconnect_2:thermocouples_sel_s1_chipselect -> thermocouples_sel:chipselect
	wire   [31:0] mm_interconnect_2_thermocouples_sel_s1_readdata;                // thermocouples_sel:readdata -> mm_interconnect_2:thermocouples_sel_s1_readdata
	wire    [1:0] mm_interconnect_2_thermocouples_sel_s1_address;                 // mm_interconnect_2:thermocouples_sel_s1_address -> thermocouples_sel:address
	wire          mm_interconnect_2_thermocouples_sel_s1_write;                   // mm_interconnect_2:thermocouples_sel_s1_write -> thermocouples_sel:write_n
	wire   [31:0] mm_interconnect_2_thermocouples_sel_s1_writedata;               // mm_interconnect_2:thermocouples_sel_s1_writedata -> thermocouples_sel:writedata
	wire          mm_interconnect_2_electrode_voltage_s1_chipselect;              // mm_interconnect_2:electrode_voltage_s1_chipselect -> electrode_voltage:chipselect
	wire   [31:0] mm_interconnect_2_electrode_voltage_s1_readdata;                // electrode_voltage:readdata -> mm_interconnect_2:electrode_voltage_s1_readdata
	wire    [1:0] mm_interconnect_2_electrode_voltage_s1_address;                 // mm_interconnect_2:electrode_voltage_s1_address -> electrode_voltage:address
	wire          mm_interconnect_2_electrode_voltage_s1_write;                   // mm_interconnect_2:electrode_voltage_s1_write -> electrode_voltage:write_n
	wire   [31:0] mm_interconnect_2_electrode_voltage_s1_writedata;               // mm_interconnect_2:electrode_voltage_s1_writedata -> electrode_voltage:writedata
	wire          mm_interconnect_2_iteration_number_s1_chipselect;               // mm_interconnect_2:iteration_number_s1_chipselect -> iteration_number:chipselect
	wire   [31:0] mm_interconnect_2_iteration_number_s1_readdata;                 // iteration_number:readdata -> mm_interconnect_2:iteration_number_s1_readdata
	wire    [1:0] mm_interconnect_2_iteration_number_s1_address;                  // mm_interconnect_2:iteration_number_s1_address -> iteration_number:address
	wire          mm_interconnect_2_iteration_number_s1_write;                    // mm_interconnect_2:iteration_number_s1_write -> iteration_number:write_n
	wire   [31:0] mm_interconnect_2_iteration_number_s1_writedata;                // mm_interconnect_2:iteration_number_s1_writedata -> iteration_number:writedata
	wire   [31:0] mm_interconnect_2_finish_fdtd_s1_readdata;                      // finish_fdtd:readdata -> mm_interconnect_2:finish_fdtd_s1_readdata
	wire    [1:0] mm_interconnect_2_finish_fdtd_s1_address;                       // mm_interconnect_2:finish_fdtd_s1_address -> finish_fdtd:address
	wire   [31:0] mm_interconnect_2_module_csr_s1_readdata;                       // module_csr:readdata -> mm_interconnect_2:module_csr_s1_readdata
	wire    [1:0] mm_interconnect_2_module_csr_s1_address;                        // mm_interconnect_2:module_csr_s1_address -> module_csr:address
	wire          mm_interconnect_2_power_unlock_s1_chipselect;                   // mm_interconnect_2:power_unlock_s1_chipselect -> power_unlock:chipselect
	wire   [31:0] mm_interconnect_2_power_unlock_s1_readdata;                     // power_unlock:readdata -> mm_interconnect_2:power_unlock_s1_readdata
	wire    [1:0] mm_interconnect_2_power_unlock_s1_address;                      // mm_interconnect_2:power_unlock_s1_address -> power_unlock:address
	wire          mm_interconnect_2_power_unlock_s1_write;                        // mm_interconnect_2:power_unlock_s1_write -> power_unlock:write_n
	wire   [31:0] mm_interconnect_2_power_unlock_s1_writedata;                    // mm_interconnect_2:power_unlock_s1_writedata -> power_unlock:writedata
	wire          mm_interconnect_2_hw_reset_s1_chipselect;                       // mm_interconnect_2:HW_reset_s1_chipselect -> HW_reset:chipselect
	wire   [31:0] mm_interconnect_2_hw_reset_s1_readdata;                         // HW_reset:readdata -> mm_interconnect_2:HW_reset_s1_readdata
	wire    [1:0] mm_interconnect_2_hw_reset_s1_address;                          // mm_interconnect_2:HW_reset_s1_address -> HW_reset:address
	wire          mm_interconnect_2_hw_reset_s1_write;                            // mm_interconnect_2:HW_reset_s1_write -> HW_reset:write_n
	wire   [31:0] mm_interconnect_2_hw_reset_s1_writedata;                        // mm_interconnect_2:HW_reset_s1_writedata -> HW_reset:writedata
	wire   [31:0] mm_interconnect_2_pixel_dma_addr_translation_slave_readdata;    // Pixel_DMA_Addr_Translation:slave_readdata -> mm_interconnect_2:Pixel_DMA_Addr_Translation_slave_readdata
	wire          mm_interconnect_2_pixel_dma_addr_translation_slave_waitrequest; // Pixel_DMA_Addr_Translation:slave_waitrequest -> mm_interconnect_2:Pixel_DMA_Addr_Translation_slave_waitrequest
	wire    [1:0] mm_interconnect_2_pixel_dma_addr_translation_slave_address;     // mm_interconnect_2:Pixel_DMA_Addr_Translation_slave_address -> Pixel_DMA_Addr_Translation:slave_address
	wire          mm_interconnect_2_pixel_dma_addr_translation_slave_read;        // mm_interconnect_2:Pixel_DMA_Addr_Translation_slave_read -> Pixel_DMA_Addr_Translation:slave_read
	wire    [3:0] mm_interconnect_2_pixel_dma_addr_translation_slave_byteenable;  // mm_interconnect_2:Pixel_DMA_Addr_Translation_slave_byteenable -> Pixel_DMA_Addr_Translation:slave_byteenable
	wire          mm_interconnect_2_pixel_dma_addr_translation_slave_write;       // mm_interconnect_2:Pixel_DMA_Addr_Translation_slave_write -> Pixel_DMA_Addr_Translation:slave_write
	wire   [31:0] mm_interconnect_2_pixel_dma_addr_translation_slave_writedata;   // mm_interconnect_2:Pixel_DMA_Addr_Translation_slave_writedata -> Pixel_DMA_Addr_Translation:slave_writedata
	wire   [31:0] pixel_dma_addr_translation_master_readdata;                     // mm_interconnect_3:Pixel_DMA_Addr_Translation_master_readdata -> Pixel_DMA_Addr_Translation:master_readdata
	wire          pixel_dma_addr_translation_master_waitrequest;                  // mm_interconnect_3:Pixel_DMA_Addr_Translation_master_waitrequest -> Pixel_DMA_Addr_Translation:master_waitrequest
	wire    [1:0] pixel_dma_addr_translation_master_address;                      // Pixel_DMA_Addr_Translation:master_address -> mm_interconnect_3:Pixel_DMA_Addr_Translation_master_address
	wire    [3:0] pixel_dma_addr_translation_master_byteenable;                   // Pixel_DMA_Addr_Translation:master_byteenable -> mm_interconnect_3:Pixel_DMA_Addr_Translation_master_byteenable
	wire          pixel_dma_addr_translation_master_read;                         // Pixel_DMA_Addr_Translation:master_read -> mm_interconnect_3:Pixel_DMA_Addr_Translation_master_read
	wire          pixel_dma_addr_translation_master_write;                        // Pixel_DMA_Addr_Translation:master_write -> mm_interconnect_3:Pixel_DMA_Addr_Translation_master_write
	wire   [31:0] pixel_dma_addr_translation_master_writedata;                    // Pixel_DMA_Addr_Translation:master_writedata -> mm_interconnect_3:Pixel_DMA_Addr_Translation_master_writedata
	wire   [31:0] mm_interconnect_3_vga_subsystem_pixel_dma_slave_readdata;       // VGA_subsystem:pixel_dma_slave_readdata -> mm_interconnect_3:VGA_subsystem_pixel_dma_slave_readdata
	wire    [1:0] mm_interconnect_3_vga_subsystem_pixel_dma_slave_address;        // mm_interconnect_3:VGA_subsystem_pixel_dma_slave_address -> VGA_subsystem:pixel_dma_slave_address
	wire          mm_interconnect_3_vga_subsystem_pixel_dma_slave_read;           // mm_interconnect_3:VGA_subsystem_pixel_dma_slave_read -> VGA_subsystem:pixel_dma_slave_read
	wire    [3:0] mm_interconnect_3_vga_subsystem_pixel_dma_slave_byteenable;     // mm_interconnect_3:VGA_subsystem_pixel_dma_slave_byteenable -> VGA_subsystem:pixel_dma_slave_byteenable
	wire          mm_interconnect_3_vga_subsystem_pixel_dma_slave_write;          // mm_interconnect_3:VGA_subsystem_pixel_dma_slave_write -> VGA_subsystem:pixel_dma_slave_write
	wire   [31:0] mm_interconnect_3_vga_subsystem_pixel_dma_slave_writedata;      // mm_interconnect_3:VGA_subsystem_pixel_dma_slave_writedata -> VGA_subsystem:pixel_dma_slave_writedata
	wire   [31:0] hps_0_f2h_irq0_irq;                                             // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                             // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [HW_reset:reset_n, Number32:reset_n, O_pw_forward:reset_n, O_pw_reversed:reset_n, O_temperature2:reset_n, O_temperature:reset_n, Pixel_DMA_Addr_Translation:reset, SP:reset_n, SW:reset_n, command_from_hps:reset_n, electrode_voltage:reset_n, fifo_FPGA_to_HPS:rdreset_n, fifo_HPS_to_FPGA:wrreset_n, finish_fdtd:reset_n, iteration_number:reset_n, mm_interconnect_1:VGA_subsystem_sys_reset_reset_bridge_in_reset_reset, mm_interconnect_1:fifo_HPS_to_FPGA_reset_in_reset_bridge_in_reset_reset, mm_interconnect_2:VGA_subsystem_sys_reset_reset_bridge_in_reset_reset, mm_interconnect_2:fifo_HPS_to_FPGA_reset_in_reset_bridge_in_reset_reset, mm_interconnect_3:Pixel_DMA_Addr_Translation_reset_reset_bridge_in_reset_reset, mm_interconnect_3:VGA_subsystem_sys_reset_reset_bridge_in_reset_reset, module_csr:reset_n, onchip_ram1:reset2, onchip_ram2:reset2, power_unlock:reset_n, rf_on_off:reset_n, rst_translator:in_reset, sdram:reset_n, thermocouples_sel:reset_n]
	wire          rst_controller_reset_out_reset_req;                             // rst_controller:reset_req -> [onchip_ram1:reset_req2, onchip_ram2:reset_req2, rst_translator:reset_req_in]
	wire          hps_0_h2f_reset_reset;                                          // hps_0:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0]
	wire          clocks_reset_source_reset;                                      // clocks:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire          rst_controller_001_reset_out_reset;                             // rst_controller_001:reset_out -> VGA_subsystem:sys_reset_reset_n
	wire          rst_controller_002_reset_out_reset;                             // rst_controller_002:reset_out -> [bridge_FPGA_tempADC:reset, mm_interconnect_0:bridge_FPGA_tempADC_reset_reset_bridge_in_reset_reset, temperature_adc:slave_reset_n]
	wire          rst_controller_003_reset_out_reset;                             // rst_controller_003:reset_out -> pll_adc:rst
	wire          rst_controller_004_reset_out_reset;                             // rst_controller_004:reset_out -> [mm_interconnect_1:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	nios2_HW_reset hw_reset (
		.clk        (clock_bridge_100_out_clk_clk),             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_2_hw_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_hw_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_hw_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_hw_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_hw_reset_s1_readdata),   //                    .readdata
		.out_port   (hw_reset_external_connection_export)       // external_connection.export
	);

	nios2_Number32 number32 (
		.clk      (clock_bridge_100_out_clk_clk),           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_2_number32_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_number32_s1_readdata), //                    .readdata
		.in_port  (number32_export)                         // external_connection.export
	);

	nios2_O_pw_forward o_pw_forward (
		.clk      (clock_bridge_100_out_clk_clk),               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_2_o_pw_forward_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_o_pw_forward_s1_readdata), //                    .readdata
		.in_port  (o_pw_forward_external_connection_export)     // external_connection.export
	);

	nios2_O_pw_forward o_pw_reversed (
		.clk      (clock_bridge_100_out_clk_clk),                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_2_o_pw_reversed_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_o_pw_reversed_s1_readdata), //                    .readdata
		.in_port  (o_pw_reversed_external_connection_export)     // external_connection.export
	);

	nios2_O_pw_forward o_temperature (
		.clk      (clock_bridge_100_out_clk_clk),                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_2_o_temperature_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_o_temperature_s1_readdata), //                    .readdata
		.in_port  (o_temperature_external_connection_export)     // external_connection.export
	);

	nios2_O_pw_forward o_temperature2 (
		.clk      (clock_bridge_100_out_clk_clk),                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_2_o_temperature2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_o_temperature2_s1_readdata), //                    .readdata
		.in_port  (o_temperature2_external_connection_export)     // external_connection.export
	);

	altera_up_avalon_video_dma_ctrl_addr_trans #(
		.ADDRESS_TRANSLATION_MASK (32'b11000000000000000000000000000000)
	) pixel_dma_addr_translation (
		.clk                (clock_bridge_100_out_clk_clk),                                   //  clock.clk
		.reset              (rst_controller_reset_out_reset),                                 //  reset.reset
		.slave_address      (mm_interconnect_2_pixel_dma_addr_translation_slave_address),     //  slave.address
		.slave_byteenable   (mm_interconnect_2_pixel_dma_addr_translation_slave_byteenable),  //       .byteenable
		.slave_read         (mm_interconnect_2_pixel_dma_addr_translation_slave_read),        //       .read
		.slave_write        (mm_interconnect_2_pixel_dma_addr_translation_slave_write),       //       .write
		.slave_writedata    (mm_interconnect_2_pixel_dma_addr_translation_slave_writedata),   //       .writedata
		.slave_readdata     (mm_interconnect_2_pixel_dma_addr_translation_slave_readdata),    //       .readdata
		.slave_waitrequest  (mm_interconnect_2_pixel_dma_addr_translation_slave_waitrequest), //       .waitrequest
		.master_readdata    (pixel_dma_addr_translation_master_readdata),                     // master.readdata
		.master_waitrequest (pixel_dma_addr_translation_master_waitrequest),                  //       .waitrequest
		.master_address     (pixel_dma_addr_translation_master_address),                      //       .address
		.master_byteenable  (pixel_dma_addr_translation_master_byteenable),                   //       .byteenable
		.master_read        (pixel_dma_addr_translation_master_read),                         //       .read
		.master_write       (pixel_dma_addr_translation_master_write),                        //       .write
		.master_writedata   (pixel_dma_addr_translation_master_writedata)                     //       .writedata
	);

	nios2_SP sp (
		.clk        (clock_bridge_100_out_clk_clk),       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_2_sp_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_sp_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_sp_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_sp_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_sp_s1_readdata),   //                    .readdata
		.out_port   (sp_external_connection_export)       // external_connection.export
	);

	nios2_SW sw (
		.clk      (clock_bridge_100_out_clk_clk),     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_2_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_sw_s1_readdata), //                    .readdata
		.in_port  (sw_external_connection_export)     // external_connection.export
	);

	nios2_VGA_subsystem vga_subsystem (
		.char_buffer_slave_byteenable   (mm_interconnect_1_vga_subsystem_char_buffer_slave_byteenable),  //   char_buffer_slave.byteenable
		.char_buffer_slave_chipselect   (mm_interconnect_1_vga_subsystem_char_buffer_slave_chipselect),  //                    .chipselect
		.char_buffer_slave_read         (mm_interconnect_1_vga_subsystem_char_buffer_slave_read),        //                    .read
		.char_buffer_slave_write        (mm_interconnect_1_vga_subsystem_char_buffer_slave_write),       //                    .write
		.char_buffer_slave_writedata    (mm_interconnect_1_vga_subsystem_char_buffer_slave_writedata),   //                    .writedata
		.char_buffer_slave_readdata     (mm_interconnect_1_vga_subsystem_char_buffer_slave_readdata),    //                    .readdata
		.char_buffer_slave_waitrequest  (mm_interconnect_1_vga_subsystem_char_buffer_slave_waitrequest), //                    .waitrequest
		.char_buffer_slave_address      (mm_interconnect_1_vga_subsystem_char_buffer_slave_address),     //                    .address
		.char_control_slave_address     (mm_interconnect_2_vga_subsystem_char_control_slave_address),    //  char_control_slave.address
		.char_control_slave_byteenable  (mm_interconnect_2_vga_subsystem_char_control_slave_byteenable), //                    .byteenable
		.char_control_slave_chipselect  (mm_interconnect_2_vga_subsystem_char_control_slave_chipselect), //                    .chipselect
		.char_control_slave_read        (mm_interconnect_2_vga_subsystem_char_control_slave_read),       //                    .read
		.char_control_slave_write       (mm_interconnect_2_vga_subsystem_char_control_slave_write),      //                    .write
		.char_control_slave_writedata   (mm_interconnect_2_vga_subsystem_char_control_slave_writedata),  //                    .writedata
		.char_control_slave_readdata    (mm_interconnect_2_vga_subsystem_char_control_slave_readdata),   //                    .readdata
		.pixel_dma_master_readdatavalid (vga_subsystem_pixel_dma_master_readdatavalid),                  //    pixel_dma_master.readdatavalid
		.pixel_dma_master_waitrequest   (vga_subsystem_pixel_dma_master_waitrequest),                    //                    .waitrequest
		.pixel_dma_master_address       (vga_subsystem_pixel_dma_master_address),                        //                    .address
		.pixel_dma_master_lock          (vga_subsystem_pixel_dma_master_lock),                           //                    .lock
		.pixel_dma_master_read          (vga_subsystem_pixel_dma_master_read),                           //                    .read
		.pixel_dma_master_readdata      (vga_subsystem_pixel_dma_master_readdata),                       //                    .readdata
		.pixel_dma_slave_address        (mm_interconnect_3_vga_subsystem_pixel_dma_slave_address),       //     pixel_dma_slave.address
		.pixel_dma_slave_byteenable     (mm_interconnect_3_vga_subsystem_pixel_dma_slave_byteenable),    //                    .byteenable
		.pixel_dma_slave_read           (mm_interconnect_3_vga_subsystem_pixel_dma_slave_read),          //                    .read
		.pixel_dma_slave_write          (mm_interconnect_3_vga_subsystem_pixel_dma_slave_write),         //                    .write
		.pixel_dma_slave_writedata      (mm_interconnect_3_vga_subsystem_pixel_dma_slave_writedata),     //                    .writedata
		.pixel_dma_slave_readdata       (mm_interconnect_3_vga_subsystem_pixel_dma_slave_readdata),      //                    .readdata
		.sys_clk_clk                    (clock_bridge_100_out_clk_clk),                                  //             sys_clk.clk
		.sys_reset_reset_n              (~rst_controller_001_reset_out_reset),                           //           sys_reset.reset_n
		.vga_out_CLK                    (vga_out_CLK),                                                   //             vga_out.CLK
		.vga_out_HS                     (vga_out_HS),                                                    //                    .HS
		.vga_out_VS                     (vga_out_VS),                                                    //                    .VS
		.vga_out_BLANK                  (vga_out_BLANK),                                                 //                    .BLANK
		.vga_out_SYNC                   (vga_out_SYNC),                                                  //                    .SYNC
		.vga_out_R                      (vga_out_R),                                                     //                    .R
		.vga_out_G                      (vga_out_G),                                                     //                    .G
		.vga_out_B                      (vga_out_B),                                                     //                    .B
		.video_pll_ref_reset_reset      (vga_ref_reset_reset),                                           // video_pll_ref_reset.reset
		.video_ref_clk_clk              (video_ref_clk_clk)                                              //       video_ref_clk.clk
	);

	nios2_bridge_FPGA_tempADC bridge_fpga_tempadc (
		.clk                (clock_bridge_0_in_clk_clk),                     //                clk.clk
		.reset              (rst_controller_002_reset_out_reset),            //              reset.reset
		.avalon_readdata    (bridge_fpga_tempadc_avalon_master_readdata),    //      avalon_master.readdata
		.avalon_waitrequest (bridge_fpga_tempadc_avalon_master_waitrequest), //                   .waitrequest
		.avalon_byteenable  (bridge_fpga_tempadc_avalon_master_byteenable),  //                   .byteenable
		.avalon_read        (bridge_fpga_tempadc_avalon_master_read),        //                   .read
		.avalon_write       (bridge_fpga_tempadc_avalon_master_write),       //                   .write
		.avalon_writedata   (bridge_fpga_tempadc_avalon_master_writedata),   //                   .writedata
		.avalon_address     (bridge_fpga_tempadc_avalon_master_address),     //                   .address
		.address            (bridge_0_external_interface_address),           // external_interface.export
		.byte_enable        (bridge_0_external_interface_byte_enable),       //                   .export
		.read               (bridge_0_external_interface_read),              //                   .export
		.write              (bridge_0_external_interface_write),             //                   .export
		.write_data         (bridge_0_external_interface_write_data),        //                   .export
		.acknowledge        (bridge_0_external_interface_acknowledge),       //                   .export
		.read_data          (bridge_0_external_interface_read_data)          //                   .export
	);

	nios2_clocks clocks (
		.ref_clk_clk        (clk_clk),                      //      ref_clk.clk
		.ref_reset_reset    (reset_reset),                  //    ref_reset.reset
		.sys_clk_clk        (clock_bridge_100_out_clk_clk), //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                //    sdram_clk.clk
		.reset_source_reset (clocks_reset_source_reset)     // reset_source.reset
	);

	nios2_command_from_hps command_from_hps (
		.clk        (clock_bridge_100_out_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_2_command_from_hps_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_command_from_hps_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_command_from_hps_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_command_from_hps_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_command_from_hps_s1_readdata),   //                    .readdata
		.out_port   (command_from_hps_external_connection_export)       // external_connection.export
	);

	nios2_command_from_hps electrode_voltage (
		.clk        (clock_bridge_100_out_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_2_electrode_voltage_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_electrode_voltage_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_electrode_voltage_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_electrode_voltage_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_electrode_voltage_s1_readdata),   //                    .readdata
		.out_port   (electrode_voltage_external_connection_export)       // external_connection.export
	);

	nios2_fifo_FPGA_to_HPS fifo_fpga_to_hps (
		.wrclock                        (fifo_fpga_to_hps_clk_in_clk),                          //    clk_in.clk
		.wrreset_n                      (fifo_fpga_to_hps_reset_in_reset_n),                    //  reset_in.reset_n
		.rdclock                        (clock_bridge_100_out_clk_clk),                         //   clk_out.clk
		.rdreset_n                      (~rst_controller_reset_out_reset),                      // reset_out.reset_n
		.avalonmm_write_slave_writedata (fifo_fpga_to_hps_in_writedata),                        //        in.writedata
		.avalonmm_write_slave_write     (fifo_fpga_to_hps_in_write),                            //          .write
		.avalonmm_read_slave_readdata   (mm_interconnect_1_fifo_fpga_to_hps_out_readdata),      //       out.readdata
		.avalonmm_read_slave_read       (mm_interconnect_1_fifo_fpga_to_hps_out_read),          //          .read
		.rdclk_control_slave_address    (mm_interconnect_2_fifo_fpga_to_hps_out_csr_address),   //   out_csr.address
		.rdclk_control_slave_read       (mm_interconnect_2_fifo_fpga_to_hps_out_csr_read),      //          .read
		.rdclk_control_slave_writedata  (mm_interconnect_2_fifo_fpga_to_hps_out_csr_writedata), //          .writedata
		.rdclk_control_slave_write      (mm_interconnect_2_fifo_fpga_to_hps_out_csr_write),     //          .write
		.rdclk_control_slave_readdata   (mm_interconnect_2_fifo_fpga_to_hps_out_csr_readdata),  //          .readdata
		.wrclk_control_slave_address    (fifo_fpga_to_hps_in_csr_address),                      //    in_csr.address
		.wrclk_control_slave_read       (fifo_fpga_to_hps_in_csr_read),                         //          .read
		.wrclk_control_slave_writedata  (fifo_fpga_to_hps_in_csr_writedata),                    //          .writedata
		.wrclk_control_slave_write      (fifo_fpga_to_hps_in_csr_write),                        //          .write
		.wrclk_control_slave_readdata   (fifo_fpga_to_hps_in_csr_readdata)                      //          .readdata
	);

	nios2_fifo_FPGA_to_HPS fifo_hps_to_fpga (
		.wrclock                        (clock_bridge_100_out_clk_clk),                        //    clk_in.clk
		.wrreset_n                      (~rst_controller_reset_out_reset),                     //  reset_in.reset_n
		.rdclock                        (fifo_hps_to_fpga_clk_out_clk),                        //   clk_out.clk
		.rdreset_n                      (fifo_hps_to_fpga_reset_out_reset_n),                  // reset_out.reset_n
		.avalonmm_write_slave_writedata (mm_interconnect_1_fifo_hps_to_fpga_in_writedata),     //        in.writedata
		.avalonmm_write_slave_write     (mm_interconnect_1_fifo_hps_to_fpga_in_write),         //          .write
		.avalonmm_read_slave_readdata   (fifo_hps_to_fpga_out_readdata),                       //       out.readdata
		.avalonmm_read_slave_read       (fifo_hps_to_fpga_out_read),                           //          .read
		.rdclk_control_slave_address    (fifo_hps_to_fpga_out_csr_address),                    //   out_csr.address
		.rdclk_control_slave_read       (fifo_hps_to_fpga_out_csr_read),                       //          .read
		.rdclk_control_slave_writedata  (fifo_hps_to_fpga_out_csr_writedata),                  //          .writedata
		.rdclk_control_slave_write      (fifo_hps_to_fpga_out_csr_write),                      //          .write
		.rdclk_control_slave_readdata   (fifo_hps_to_fpga_out_csr_readdata),                   //          .readdata
		.wrclk_control_slave_address    (mm_interconnect_2_fifo_hps_to_fpga_in_csr_address),   //    in_csr.address
		.wrclk_control_slave_read       (mm_interconnect_2_fifo_hps_to_fpga_in_csr_read),      //          .read
		.wrclk_control_slave_writedata  (mm_interconnect_2_fifo_hps_to_fpga_in_csr_writedata), //          .writedata
		.wrclk_control_slave_write      (mm_interconnect_2_fifo_hps_to_fpga_in_csr_write),     //          .write
		.wrclk_control_slave_readdata   (mm_interconnect_2_fifo_hps_to_fpga_in_csr_readdata)   //          .readdata
	);

	nios2_finish_fdtd finish_fdtd (
		.clk      (clock_bridge_100_out_clk_clk),              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_2_finish_fdtd_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_finish_fdtd_s1_readdata), //                    .readdata
		.in_port  (finish_fdtd_external_connection_export)     // external_connection.export
	);

	nios2_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (3)
	) hps_0 (
		.mem_a                    (memory_mem_a),                    //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                   //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                   //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                 //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                  //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                 //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                 //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),              //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                   //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                  //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                  //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                   //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK), //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL), //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL), //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK), //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),   //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),     //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),     //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),     //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),     //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),     //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),     //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),     //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),    //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),   //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),   //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),    //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),     //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),     //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),     //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),     //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),     //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),  //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),  //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),  //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),  //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),  //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),  //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk              (clock_bridge_100_out_clk_clk),    //     h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),       //    h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),     //                  .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),      //                  .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),     //                  .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),    //                  .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),     //                  .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),    //                  .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),     //                  .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),    //                  .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),    //                  .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),        //                  .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),      //                  .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),      //                  .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),      //                  .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),     //                  .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),     //                  .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),        //                  .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),      //                  .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),     //                  .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),     //                  .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),       //                  .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),     //                  .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),      //                  .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),     //                  .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),    //                  .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),     //                  .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),    //                  .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),     //                  .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),    //                  .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),    //                  .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),        //                  .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),      //                  .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),      //                  .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),      //                  .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),     //                  .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),     //                  .rready
		.f2h_axi_clk              (clock_bridge_100_out_clk_clk),    //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                //                  .awaddr
		.f2h_AWLEN                (),                                //                  .awlen
		.f2h_AWSIZE               (),                                //                  .awsize
		.f2h_AWBURST              (),                                //                  .awburst
		.f2h_AWLOCK               (),                                //                  .awlock
		.f2h_AWCACHE              (),                                //                  .awcache
		.f2h_AWPROT               (),                                //                  .awprot
		.f2h_AWVALID              (),                                //                  .awvalid
		.f2h_AWREADY              (),                                //                  .awready
		.f2h_AWUSER               (),                                //                  .awuser
		.f2h_WID                  (),                                //                  .wid
		.f2h_WDATA                (),                                //                  .wdata
		.f2h_WSTRB                (),                                //                  .wstrb
		.f2h_WLAST                (),                                //                  .wlast
		.f2h_WVALID               (),                                //                  .wvalid
		.f2h_WREADY               (),                                //                  .wready
		.f2h_BID                  (),                                //                  .bid
		.f2h_BRESP                (),                                //                  .bresp
		.f2h_BVALID               (),                                //                  .bvalid
		.f2h_BREADY               (),                                //                  .bready
		.f2h_ARID                 (),                                //                  .arid
		.f2h_ARADDR               (),                                //                  .araddr
		.f2h_ARLEN                (),                                //                  .arlen
		.f2h_ARSIZE               (),                                //                  .arsize
		.f2h_ARBURST              (),                                //                  .arburst
		.f2h_ARLOCK               (),                                //                  .arlock
		.f2h_ARCACHE              (),                                //                  .arcache
		.f2h_ARPROT               (),                                //                  .arprot
		.f2h_ARVALID              (),                                //                  .arvalid
		.f2h_ARREADY              (),                                //                  .arready
		.f2h_ARUSER               (),                                //                  .aruser
		.f2h_RID                  (),                                //                  .rid
		.f2h_RDATA                (),                                //                  .rdata
		.f2h_RRESP                (),                                //                  .rresp
		.f2h_RLAST                (),                                //                  .rlast
		.f2h_RVALID               (),                                //                  .rvalid
		.f2h_RREADY               (),                                //                  .rready
		.h2f_lw_axi_clk           (clock_bridge_100_out_clk_clk),    //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),  //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),              //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)               //          f2h_irq1.irq
	);

	nios2_iteration_number iteration_number (
		.clk        (clock_bridge_100_out_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_2_iteration_number_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_iteration_number_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_iteration_number_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_iteration_number_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_iteration_number_s1_readdata),   //                    .readdata
		.out_port   (iteration_number_external_connection_export)       // external_connection.export
	);

	nios2_O_pw_forward module_csr (
		.clk      (clock_bridge_100_out_clk_clk),             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_2_module_csr_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_module_csr_s1_readdata), //                    .readdata
		.in_port  (module_csr_external_connection_export)     // external_connection.export
	);

	nios2_onchip_ram1 onchip_ram1 (
		.clk         (clock_bridge_65_out_clk_clk),                 //   clk1.clk
		.address     (onchip_ram1_s1_address),                      //     s1.address
		.clken       (onchip_ram1_s1_clken),                        //       .clken
		.chipselect  (onchip_ram1_s1_chipselect),                   //       .chipselect
		.write       (onchip_ram1_s1_write),                        //       .write
		.readdata    (onchip_ram1_s1_readdata),                     //       .readdata
		.writedata   (onchip_ram1_s1_writedata),                    //       .writedata
		.byteenable  (onchip_ram1_s1_byteenable),                   //       .byteenable
		.reset       (onchip_ram1_reset1_reset),                    // reset1.reset
		.reset_req   (onchip_ram1_reset1_reset_req),                //       .reset_req
		.address2    (mm_interconnect_1_onchip_ram1_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_1_onchip_ram1_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_1_onchip_ram1_s2_clken),      //       .clken
		.write2      (mm_interconnect_1_onchip_ram1_s2_write),      //       .write
		.readdata2   (mm_interconnect_1_onchip_ram1_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_1_onchip_ram1_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_1_onchip_ram1_s2_byteenable), //       .byteenable
		.clk2        (clock_bridge_100_out_clk_clk),                //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),              // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	nios2_onchip_ram2 onchip_ram2 (
		.clk         (clock_bridge_65_out_clk_clk),                 //   clk1.clk
		.address     (onchip_ram2_s1_address),                      //     s1.address
		.clken       (onchip_ram2_s1_clken),                        //       .clken
		.chipselect  (onchip_ram2_s1_chipselect),                   //       .chipselect
		.write       (onchip_ram2_s1_write),                        //       .write
		.readdata    (onchip_ram2_s1_readdata),                     //       .readdata
		.writedata   (onchip_ram2_s1_writedata),                    //       .writedata
		.byteenable  (onchip_ram2_s1_byteenable),                   //       .byteenable
		.reset       (onchip_ram2_reset1_reset),                    // reset1.reset
		.reset_req   (onchip_ram2_reset1_reset_req),                //       .reset_req
		.address2    (mm_interconnect_1_onchip_ram2_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_1_onchip_ram2_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_1_onchip_ram2_s2_clken),      //       .clken
		.write2      (mm_interconnect_1_onchip_ram2_s2_write),      //       .write
		.readdata2   (mm_interconnect_1_onchip_ram2_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_1_onchip_ram2_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_1_onchip_ram2_s2_byteenable), //       .byteenable
		.clk2        (clock_bridge_100_out_clk_clk),                //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),              // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	nios2_pll_adc pll_adc (
		.refclk   (clock_bridge_100_out_clk_clk),       //  refclk.clk
		.rst      (rst_controller_003_reset_out_reset), //   reset.reset
		.outclk_0 (pll_adc_outclk0_clk),                // outclk0.clk
		.outclk_1 (clock_bridge_65_out_clk_clk),        // outclk1.clk
		.locked   (pll_adc_locked_export)               //  locked.export
	);

	nios2_HW_reset power_unlock (
		.clk        (clock_bridge_100_out_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_2_power_unlock_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_power_unlock_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_power_unlock_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_power_unlock_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_power_unlock_s1_readdata),   //                    .readdata
		.out_port   (power_unlock_external_connection_export)       // external_connection.export
	);

	nios2_rf_on_off rf_on_off (
		.clk        (clock_bridge_100_out_clk_clk),              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_2_rf_on_off_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_rf_on_off_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_rf_on_off_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_rf_on_off_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_rf_on_off_s1_readdata),   //                    .readdata
		.out_port   (rf_on_off_external_connection_export)       // external_connection.export
	);

	nios2_sdram sdram (
		.clk            (clock_bridge_100_out_clk_clk),             //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_1_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	adc_ltc2308_fifo temperature_adc (
		.slave_chipselect_n (~mm_interconnect_0_temperature_adc_slave_chipselect), //          slave.chipselect_n
		.slave_read_n       (~mm_interconnect_0_temperature_adc_slave_read),       //               .read_n
		.slave_readdata     (mm_interconnect_0_temperature_adc_slave_readdata),    //               .readdata
		.slave_addr         (mm_interconnect_0_temperature_adc_slave_address),     //               .address
		.slave_wrtie_n      (~mm_interconnect_0_temperature_adc_slave_write),      //               .write_n
		.slave_wriredata    (mm_interconnect_0_temperature_adc_slave_writedata),   //               .writedata
		.ADC_CONVST         (adc_ltc2308_0_conduit_end_CONVST),                    //    conduit_end.export
		.ADC_SCK            (adc_ltc2308_0_conduit_end_SCK),                       //               .export
		.ADC_SDI            (adc_ltc2308_0_conduit_end_SDI),                       //               .export
		.ADC_SDO            (adc_ltc2308_0_conduit_end_SDO),                       //               .export
		.slave_reset_n      (~rst_controller_002_reset_out_reset),                 //     reset_sink.reset_n
		.slave_clk          (clock_bridge_0_in_clk_clk),                           //     clock_sink.clk
		.adc_clk            (pll_adc_outclk0_clk)                                  // clock_sink_adc.clk
	);

	nios2_rf_on_off thermocouples_sel (
		.clk        (clock_bridge_100_out_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_2_thermocouples_sel_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_thermocouples_sel_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_thermocouples_sel_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_thermocouples_sel_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_thermocouples_sel_s1_readdata),   //                    .readdata
		.out_port   (thermocouples_sel_external_connection_export)       // external_connection.export
	);

	nios2_mm_interconnect_0 mm_interconnect_0 (
		.clock_bridge_0_out_clk_clk                            (clock_bridge_0_in_clk_clk),                          //                          clock_bridge_0_out_clk.clk
		.bridge_FPGA_tempADC_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                 // bridge_FPGA_tempADC_reset_reset_bridge_in_reset.reset
		.bridge_FPGA_tempADC_avalon_master_address             (bridge_fpga_tempadc_avalon_master_address),          //               bridge_FPGA_tempADC_avalon_master.address
		.bridge_FPGA_tempADC_avalon_master_waitrequest         (bridge_fpga_tempadc_avalon_master_waitrequest),      //                                                .waitrequest
		.bridge_FPGA_tempADC_avalon_master_byteenable          (bridge_fpga_tempadc_avalon_master_byteenable),       //                                                .byteenable
		.bridge_FPGA_tempADC_avalon_master_read                (bridge_fpga_tempadc_avalon_master_read),             //                                                .read
		.bridge_FPGA_tempADC_avalon_master_readdata            (bridge_fpga_tempadc_avalon_master_readdata),         //                                                .readdata
		.bridge_FPGA_tempADC_avalon_master_write               (bridge_fpga_tempadc_avalon_master_write),            //                                                .write
		.bridge_FPGA_tempADC_avalon_master_writedata           (bridge_fpga_tempadc_avalon_master_writedata),        //                                                .writedata
		.temperature_adc_slave_address                         (mm_interconnect_0_temperature_adc_slave_address),    //                           temperature_adc_slave.address
		.temperature_adc_slave_write                           (mm_interconnect_0_temperature_adc_slave_write),      //                                                .write
		.temperature_adc_slave_read                            (mm_interconnect_0_temperature_adc_slave_read),       //                                                .read
		.temperature_adc_slave_readdata                        (mm_interconnect_0_temperature_adc_slave_readdata),   //                                                .readdata
		.temperature_adc_slave_writedata                       (mm_interconnect_0_temperature_adc_slave_writedata),  //                                                .writedata
		.temperature_adc_slave_chipselect                      (mm_interconnect_0_temperature_adc_slave_chipselect)  //                                                .chipselect
	);

	nios2_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                                     //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                                   //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                                    //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                                   //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                                  //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                                   //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                                  //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                                   //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                                  //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                                  //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                                      //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                                    //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                                    //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                                    //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                                   //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                                   //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                                      //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                                    //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                                   //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                                   //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                                     //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                                   //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                                    //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                                   //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                                  //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                                   //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                                  //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                                   //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                                  //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                                  //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                                      //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                                    //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                                    //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                                    //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                                   //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                                   //                                                           .rready
		.clocks_sys_clk_clk                                               (clock_bridge_100_out_clk_clk),                                  //                                             clocks_sys_clk.clk
		.fifo_HPS_to_FPGA_reset_in_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                                //            fifo_HPS_to_FPGA_reset_in_reset_bridge_in_reset.reset
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                            // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.VGA_subsystem_sys_reset_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                                //              VGA_subsystem_sys_reset_reset_bridge_in_reset.reset
		.VGA_subsystem_pixel_dma_master_address                           (vga_subsystem_pixel_dma_master_address),                        //                             VGA_subsystem_pixel_dma_master.address
		.VGA_subsystem_pixel_dma_master_waitrequest                       (vga_subsystem_pixel_dma_master_waitrequest),                    //                                                           .waitrequest
		.VGA_subsystem_pixel_dma_master_read                              (vga_subsystem_pixel_dma_master_read),                           //                                                           .read
		.VGA_subsystem_pixel_dma_master_readdata                          (vga_subsystem_pixel_dma_master_readdata),                       //                                                           .readdata
		.VGA_subsystem_pixel_dma_master_readdatavalid                     (vga_subsystem_pixel_dma_master_readdatavalid),                  //                                                           .readdatavalid
		.VGA_subsystem_pixel_dma_master_lock                              (vga_subsystem_pixel_dma_master_lock),                           //                                                           .lock
		.fifo_FPGA_to_HPS_out_read                                        (mm_interconnect_1_fifo_fpga_to_hps_out_read),                   //                                       fifo_FPGA_to_HPS_out.read
		.fifo_FPGA_to_HPS_out_readdata                                    (mm_interconnect_1_fifo_fpga_to_hps_out_readdata),               //                                                           .readdata
		.fifo_HPS_to_FPGA_in_write                                        (mm_interconnect_1_fifo_hps_to_fpga_in_write),                   //                                        fifo_HPS_to_FPGA_in.write
		.fifo_HPS_to_FPGA_in_writedata                                    (mm_interconnect_1_fifo_hps_to_fpga_in_writedata),               //                                                           .writedata
		.onchip_ram1_s2_address                                           (mm_interconnect_1_onchip_ram1_s2_address),                      //                                             onchip_ram1_s2.address
		.onchip_ram1_s2_write                                             (mm_interconnect_1_onchip_ram1_s2_write),                        //                                                           .write
		.onchip_ram1_s2_readdata                                          (mm_interconnect_1_onchip_ram1_s2_readdata),                     //                                                           .readdata
		.onchip_ram1_s2_writedata                                         (mm_interconnect_1_onchip_ram1_s2_writedata),                    //                                                           .writedata
		.onchip_ram1_s2_byteenable                                        (mm_interconnect_1_onchip_ram1_s2_byteenable),                   //                                                           .byteenable
		.onchip_ram1_s2_chipselect                                        (mm_interconnect_1_onchip_ram1_s2_chipselect),                   //                                                           .chipselect
		.onchip_ram1_s2_clken                                             (mm_interconnect_1_onchip_ram1_s2_clken),                        //                                                           .clken
		.onchip_ram2_s2_address                                           (mm_interconnect_1_onchip_ram2_s2_address),                      //                                             onchip_ram2_s2.address
		.onchip_ram2_s2_write                                             (mm_interconnect_1_onchip_ram2_s2_write),                        //                                                           .write
		.onchip_ram2_s2_readdata                                          (mm_interconnect_1_onchip_ram2_s2_readdata),                     //                                                           .readdata
		.onchip_ram2_s2_writedata                                         (mm_interconnect_1_onchip_ram2_s2_writedata),                    //                                                           .writedata
		.onchip_ram2_s2_byteenable                                        (mm_interconnect_1_onchip_ram2_s2_byteenable),                   //                                                           .byteenable
		.onchip_ram2_s2_chipselect                                        (mm_interconnect_1_onchip_ram2_s2_chipselect),                   //                                                           .chipselect
		.onchip_ram2_s2_clken                                             (mm_interconnect_1_onchip_ram2_s2_clken),                        //                                                           .clken
		.sdram_s1_address                                                 (mm_interconnect_1_sdram_s1_address),                            //                                                   sdram_s1.address
		.sdram_s1_write                                                   (mm_interconnect_1_sdram_s1_write),                              //                                                           .write
		.sdram_s1_read                                                    (mm_interconnect_1_sdram_s1_read),                               //                                                           .read
		.sdram_s1_readdata                                                (mm_interconnect_1_sdram_s1_readdata),                           //                                                           .readdata
		.sdram_s1_writedata                                               (mm_interconnect_1_sdram_s1_writedata),                          //                                                           .writedata
		.sdram_s1_byteenable                                              (mm_interconnect_1_sdram_s1_byteenable),                         //                                                           .byteenable
		.sdram_s1_readdatavalid                                           (mm_interconnect_1_sdram_s1_readdatavalid),                      //                                                           .readdatavalid
		.sdram_s1_waitrequest                                             (mm_interconnect_1_sdram_s1_waitrequest),                        //                                                           .waitrequest
		.sdram_s1_chipselect                                              (mm_interconnect_1_sdram_s1_chipselect),                         //                                                           .chipselect
		.VGA_subsystem_char_buffer_slave_address                          (mm_interconnect_1_vga_subsystem_char_buffer_slave_address),     //                            VGA_subsystem_char_buffer_slave.address
		.VGA_subsystem_char_buffer_slave_write                            (mm_interconnect_1_vga_subsystem_char_buffer_slave_write),       //                                                           .write
		.VGA_subsystem_char_buffer_slave_read                             (mm_interconnect_1_vga_subsystem_char_buffer_slave_read),        //                                                           .read
		.VGA_subsystem_char_buffer_slave_readdata                         (mm_interconnect_1_vga_subsystem_char_buffer_slave_readdata),    //                                                           .readdata
		.VGA_subsystem_char_buffer_slave_writedata                        (mm_interconnect_1_vga_subsystem_char_buffer_slave_writedata),   //                                                           .writedata
		.VGA_subsystem_char_buffer_slave_byteenable                       (mm_interconnect_1_vga_subsystem_char_buffer_slave_byteenable),  //                                                           .byteenable
		.VGA_subsystem_char_buffer_slave_waitrequest                      (mm_interconnect_1_vga_subsystem_char_buffer_slave_waitrequest), //                                                           .waitrequest
		.VGA_subsystem_char_buffer_slave_chipselect                       (mm_interconnect_1_vga_subsystem_char_buffer_slave_chipselect)   //                                                           .chipselect
	);

	nios2_mm_interconnect_2 mm_interconnect_2 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                   //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                                 //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                                  //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                                 //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                                //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                                 //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                                //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                                 //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                                //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                                //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                    //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                                  //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                                  //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                                  //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                                 //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                                 //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                    //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                                  //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                                 //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                                 //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                   //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                                 //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                                  //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                                 //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                                //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                                 //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                                //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                                 //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                                //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                                //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                    //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                                  //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                                  //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                                  //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                                 //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                                 //                                                              .rready
		.clocks_sys_clk_clk                                                  (clock_bridge_100_out_clk_clk),                                   //                                                clocks_sys_clk.clk
		.fifo_HPS_to_FPGA_reset_in_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                                 //               fifo_HPS_to_FPGA_reset_in_reset_bridge_in_reset.reset
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                             // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.VGA_subsystem_sys_reset_reset_bridge_in_reset_reset                 (rst_controller_reset_out_reset),                                 //                 VGA_subsystem_sys_reset_reset_bridge_in_reset.reset
		.command_from_hps_s1_address                                         (mm_interconnect_2_command_from_hps_s1_address),                  //                                           command_from_hps_s1.address
		.command_from_hps_s1_write                                           (mm_interconnect_2_command_from_hps_s1_write),                    //                                                              .write
		.command_from_hps_s1_readdata                                        (mm_interconnect_2_command_from_hps_s1_readdata),                 //                                                              .readdata
		.command_from_hps_s1_writedata                                       (mm_interconnect_2_command_from_hps_s1_writedata),                //                                                              .writedata
		.command_from_hps_s1_chipselect                                      (mm_interconnect_2_command_from_hps_s1_chipselect),               //                                                              .chipselect
		.electrode_voltage_s1_address                                        (mm_interconnect_2_electrode_voltage_s1_address),                 //                                          electrode_voltage_s1.address
		.electrode_voltage_s1_write                                          (mm_interconnect_2_electrode_voltage_s1_write),                   //                                                              .write
		.electrode_voltage_s1_readdata                                       (mm_interconnect_2_electrode_voltage_s1_readdata),                //                                                              .readdata
		.electrode_voltage_s1_writedata                                      (mm_interconnect_2_electrode_voltage_s1_writedata),               //                                                              .writedata
		.electrode_voltage_s1_chipselect                                     (mm_interconnect_2_electrode_voltage_s1_chipselect),              //                                                              .chipselect
		.fifo_FPGA_to_HPS_out_csr_address                                    (mm_interconnect_2_fifo_fpga_to_hps_out_csr_address),             //                                      fifo_FPGA_to_HPS_out_csr.address
		.fifo_FPGA_to_HPS_out_csr_write                                      (mm_interconnect_2_fifo_fpga_to_hps_out_csr_write),               //                                                              .write
		.fifo_FPGA_to_HPS_out_csr_read                                       (mm_interconnect_2_fifo_fpga_to_hps_out_csr_read),                //                                                              .read
		.fifo_FPGA_to_HPS_out_csr_readdata                                   (mm_interconnect_2_fifo_fpga_to_hps_out_csr_readdata),            //                                                              .readdata
		.fifo_FPGA_to_HPS_out_csr_writedata                                  (mm_interconnect_2_fifo_fpga_to_hps_out_csr_writedata),           //                                                              .writedata
		.fifo_HPS_to_FPGA_in_csr_address                                     (mm_interconnect_2_fifo_hps_to_fpga_in_csr_address),              //                                       fifo_HPS_to_FPGA_in_csr.address
		.fifo_HPS_to_FPGA_in_csr_write                                       (mm_interconnect_2_fifo_hps_to_fpga_in_csr_write),                //                                                              .write
		.fifo_HPS_to_FPGA_in_csr_read                                        (mm_interconnect_2_fifo_hps_to_fpga_in_csr_read),                 //                                                              .read
		.fifo_HPS_to_FPGA_in_csr_readdata                                    (mm_interconnect_2_fifo_hps_to_fpga_in_csr_readdata),             //                                                              .readdata
		.fifo_HPS_to_FPGA_in_csr_writedata                                   (mm_interconnect_2_fifo_hps_to_fpga_in_csr_writedata),            //                                                              .writedata
		.finish_fdtd_s1_address                                              (mm_interconnect_2_finish_fdtd_s1_address),                       //                                                finish_fdtd_s1.address
		.finish_fdtd_s1_readdata                                             (mm_interconnect_2_finish_fdtd_s1_readdata),                      //                                                              .readdata
		.HW_reset_s1_address                                                 (mm_interconnect_2_hw_reset_s1_address),                          //                                                   HW_reset_s1.address
		.HW_reset_s1_write                                                   (mm_interconnect_2_hw_reset_s1_write),                            //                                                              .write
		.HW_reset_s1_readdata                                                (mm_interconnect_2_hw_reset_s1_readdata),                         //                                                              .readdata
		.HW_reset_s1_writedata                                               (mm_interconnect_2_hw_reset_s1_writedata),                        //                                                              .writedata
		.HW_reset_s1_chipselect                                              (mm_interconnect_2_hw_reset_s1_chipselect),                       //                                                              .chipselect
		.iteration_number_s1_address                                         (mm_interconnect_2_iteration_number_s1_address),                  //                                           iteration_number_s1.address
		.iteration_number_s1_write                                           (mm_interconnect_2_iteration_number_s1_write),                    //                                                              .write
		.iteration_number_s1_readdata                                        (mm_interconnect_2_iteration_number_s1_readdata),                 //                                                              .readdata
		.iteration_number_s1_writedata                                       (mm_interconnect_2_iteration_number_s1_writedata),                //                                                              .writedata
		.iteration_number_s1_chipselect                                      (mm_interconnect_2_iteration_number_s1_chipselect),               //                                                              .chipselect
		.module_csr_s1_address                                               (mm_interconnect_2_module_csr_s1_address),                        //                                                 module_csr_s1.address
		.module_csr_s1_readdata                                              (mm_interconnect_2_module_csr_s1_readdata),                       //                                                              .readdata
		.Number32_s1_address                                                 (mm_interconnect_2_number32_s1_address),                          //                                                   Number32_s1.address
		.Number32_s1_readdata                                                (mm_interconnect_2_number32_s1_readdata),                         //                                                              .readdata
		.O_pw_forward_s1_address                                             (mm_interconnect_2_o_pw_forward_s1_address),                      //                                               O_pw_forward_s1.address
		.O_pw_forward_s1_readdata                                            (mm_interconnect_2_o_pw_forward_s1_readdata),                     //                                                              .readdata
		.O_pw_reversed_s1_address                                            (mm_interconnect_2_o_pw_reversed_s1_address),                     //                                              O_pw_reversed_s1.address
		.O_pw_reversed_s1_readdata                                           (mm_interconnect_2_o_pw_reversed_s1_readdata),                    //                                                              .readdata
		.O_temperature_s1_address                                            (mm_interconnect_2_o_temperature_s1_address),                     //                                              O_temperature_s1.address
		.O_temperature_s1_readdata                                           (mm_interconnect_2_o_temperature_s1_readdata),                    //                                                              .readdata
		.O_temperature2_s1_address                                           (mm_interconnect_2_o_temperature2_s1_address),                    //                                             O_temperature2_s1.address
		.O_temperature2_s1_readdata                                          (mm_interconnect_2_o_temperature2_s1_readdata),                   //                                                              .readdata
		.Pixel_DMA_Addr_Translation_slave_address                            (mm_interconnect_2_pixel_dma_addr_translation_slave_address),     //                              Pixel_DMA_Addr_Translation_slave.address
		.Pixel_DMA_Addr_Translation_slave_write                              (mm_interconnect_2_pixel_dma_addr_translation_slave_write),       //                                                              .write
		.Pixel_DMA_Addr_Translation_slave_read                               (mm_interconnect_2_pixel_dma_addr_translation_slave_read),        //                                                              .read
		.Pixel_DMA_Addr_Translation_slave_readdata                           (mm_interconnect_2_pixel_dma_addr_translation_slave_readdata),    //                                                              .readdata
		.Pixel_DMA_Addr_Translation_slave_writedata                          (mm_interconnect_2_pixel_dma_addr_translation_slave_writedata),   //                                                              .writedata
		.Pixel_DMA_Addr_Translation_slave_byteenable                         (mm_interconnect_2_pixel_dma_addr_translation_slave_byteenable),  //                                                              .byteenable
		.Pixel_DMA_Addr_Translation_slave_waitrequest                        (mm_interconnect_2_pixel_dma_addr_translation_slave_waitrequest), //                                                              .waitrequest
		.power_unlock_s1_address                                             (mm_interconnect_2_power_unlock_s1_address),                      //                                               power_unlock_s1.address
		.power_unlock_s1_write                                               (mm_interconnect_2_power_unlock_s1_write),                        //                                                              .write
		.power_unlock_s1_readdata                                            (mm_interconnect_2_power_unlock_s1_readdata),                     //                                                              .readdata
		.power_unlock_s1_writedata                                           (mm_interconnect_2_power_unlock_s1_writedata),                    //                                                              .writedata
		.power_unlock_s1_chipselect                                          (mm_interconnect_2_power_unlock_s1_chipselect),                   //                                                              .chipselect
		.rf_on_off_s1_address                                                (mm_interconnect_2_rf_on_off_s1_address),                         //                                                  rf_on_off_s1.address
		.rf_on_off_s1_write                                                  (mm_interconnect_2_rf_on_off_s1_write),                           //                                                              .write
		.rf_on_off_s1_readdata                                               (mm_interconnect_2_rf_on_off_s1_readdata),                        //                                                              .readdata
		.rf_on_off_s1_writedata                                              (mm_interconnect_2_rf_on_off_s1_writedata),                       //                                                              .writedata
		.rf_on_off_s1_chipselect                                             (mm_interconnect_2_rf_on_off_s1_chipselect),                      //                                                              .chipselect
		.SP_s1_address                                                       (mm_interconnect_2_sp_s1_address),                                //                                                         SP_s1.address
		.SP_s1_write                                                         (mm_interconnect_2_sp_s1_write),                                  //                                                              .write
		.SP_s1_readdata                                                      (mm_interconnect_2_sp_s1_readdata),                               //                                                              .readdata
		.SP_s1_writedata                                                     (mm_interconnect_2_sp_s1_writedata),                              //                                                              .writedata
		.SP_s1_chipselect                                                    (mm_interconnect_2_sp_s1_chipselect),                             //                                                              .chipselect
		.SW_s1_address                                                       (mm_interconnect_2_sw_s1_address),                                //                                                         SW_s1.address
		.SW_s1_readdata                                                      (mm_interconnect_2_sw_s1_readdata),                               //                                                              .readdata
		.thermocouples_sel_s1_address                                        (mm_interconnect_2_thermocouples_sel_s1_address),                 //                                          thermocouples_sel_s1.address
		.thermocouples_sel_s1_write                                          (mm_interconnect_2_thermocouples_sel_s1_write),                   //                                                              .write
		.thermocouples_sel_s1_readdata                                       (mm_interconnect_2_thermocouples_sel_s1_readdata),                //                                                              .readdata
		.thermocouples_sel_s1_writedata                                      (mm_interconnect_2_thermocouples_sel_s1_writedata),               //                                                              .writedata
		.thermocouples_sel_s1_chipselect                                     (mm_interconnect_2_thermocouples_sel_s1_chipselect),              //                                                              .chipselect
		.VGA_subsystem_char_control_slave_address                            (mm_interconnect_2_vga_subsystem_char_control_slave_address),     //                              VGA_subsystem_char_control_slave.address
		.VGA_subsystem_char_control_slave_write                              (mm_interconnect_2_vga_subsystem_char_control_slave_write),       //                                                              .write
		.VGA_subsystem_char_control_slave_read                               (mm_interconnect_2_vga_subsystem_char_control_slave_read),        //                                                              .read
		.VGA_subsystem_char_control_slave_readdata                           (mm_interconnect_2_vga_subsystem_char_control_slave_readdata),    //                                                              .readdata
		.VGA_subsystem_char_control_slave_writedata                          (mm_interconnect_2_vga_subsystem_char_control_slave_writedata),   //                                                              .writedata
		.VGA_subsystem_char_control_slave_byteenable                         (mm_interconnect_2_vga_subsystem_char_control_slave_byteenable),  //                                                              .byteenable
		.VGA_subsystem_char_control_slave_chipselect                         (mm_interconnect_2_vga_subsystem_char_control_slave_chipselect)   //                                                              .chipselect
	);

	nios2_mm_interconnect_3 mm_interconnect_3 (
		.clocks_sys_clk_clk                                           (clock_bridge_100_out_clk_clk),                               //                                         clocks_sys_clk.clk
		.Pixel_DMA_Addr_Translation_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // Pixel_DMA_Addr_Translation_reset_reset_bridge_in_reset.reset
		.VGA_subsystem_sys_reset_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                             //          VGA_subsystem_sys_reset_reset_bridge_in_reset.reset
		.Pixel_DMA_Addr_Translation_master_address                    (pixel_dma_addr_translation_master_address),                  //                      Pixel_DMA_Addr_Translation_master.address
		.Pixel_DMA_Addr_Translation_master_waitrequest                (pixel_dma_addr_translation_master_waitrequest),              //                                                       .waitrequest
		.Pixel_DMA_Addr_Translation_master_byteenable                 (pixel_dma_addr_translation_master_byteenable),               //                                                       .byteenable
		.Pixel_DMA_Addr_Translation_master_read                       (pixel_dma_addr_translation_master_read),                     //                                                       .read
		.Pixel_DMA_Addr_Translation_master_readdata                   (pixel_dma_addr_translation_master_readdata),                 //                                                       .readdata
		.Pixel_DMA_Addr_Translation_master_write                      (pixel_dma_addr_translation_master_write),                    //                                                       .write
		.Pixel_DMA_Addr_Translation_master_writedata                  (pixel_dma_addr_translation_master_writedata),                //                                                       .writedata
		.VGA_subsystem_pixel_dma_slave_address                        (mm_interconnect_3_vga_subsystem_pixel_dma_slave_address),    //                          VGA_subsystem_pixel_dma_slave.address
		.VGA_subsystem_pixel_dma_slave_write                          (mm_interconnect_3_vga_subsystem_pixel_dma_slave_write),      //                                                       .write
		.VGA_subsystem_pixel_dma_slave_read                           (mm_interconnect_3_vga_subsystem_pixel_dma_slave_read),       //                                                       .read
		.VGA_subsystem_pixel_dma_slave_readdata                       (mm_interconnect_3_vga_subsystem_pixel_dma_slave_readdata),   //                                                       .readdata
		.VGA_subsystem_pixel_dma_slave_writedata                      (mm_interconnect_3_vga_subsystem_pixel_dma_slave_writedata),  //                                                       .writedata
		.VGA_subsystem_pixel_dma_slave_byteenable                     (mm_interconnect_3_vga_subsystem_pixel_dma_slave_byteenable)  //                                                       .byteenable
	);

	nios2_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	nios2_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.reset_in1      (clocks_reset_source_reset),          // reset_in1.reset
		.clk            (clock_bridge_100_out_clk_clk),       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.reset_in1      (clocks_reset_source_reset),          // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.reset_in1      (clocks_reset_source_reset),          // reset_in1.reset
		.clk            (clock_bridge_0_in_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.reset_in1      (clocks_reset_source_reset),          // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clock_bridge_100_out_clk_clk),       //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
